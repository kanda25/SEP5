module sevenSeg(
  input [3:0] D;
  output [6:0] Q;
);

always @(D);
  

endmodule