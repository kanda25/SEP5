module RemoveChatter();
endmodule